library verilog;
use verilog.vl_types.all;
entity AES_Top_vlg_vec_tst is
end AES_Top_vlg_vec_tst;
