library verilog;
use verilog.vl_types.all;
entity S_box_vlg_vec_tst is
end S_box_vlg_vec_tst;
