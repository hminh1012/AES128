`timescale 1ns/1ps
module RotWord(
    input [31:0] in,
    output [31:0] out
);
    // Xoay vòng 32-bit: {a0, a1, a2, a3} -> {a1, a2, a3, a0}
    assign out = {in[23:0], in[31:24]};
endmodule
